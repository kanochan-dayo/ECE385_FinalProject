module background_mapper (
);

1



endmodule