module key_f(input [7:0] addr, 
output [15:0] key_1, 
output [15:0] key_2, 
output [15:0] key_3, 
output [15:0] key_4);
parameter [0:255][15:0] mem={
16'b0000000001000111,        // LineF00 1.199at index 3
16'b0000000001111101,        // LineF00 2.099at index 6
16'b0000000010110010,        // LineF00 2.998at index 8
16'b0000000011000110,        // LineF00 3.332at index 10
16'b0000000110000011,        // LineF00 6.499at index 18
16'b0000000110010111,        // LineF00 6.831at index 20
16'b0000000110111000,        // LineF00 7.399at index 22
16'b0000001000000000,        // LineF00 8.598at index 25
16'b0000001001000001,        // LineF00 9.700at index 28
16'b0100001001101011,        // LineF01 10.398at index 30
16'b1000001101010011,        // LineF10 14.298at index 33
16'b0000001110111010,        // LineF00 16.033at index 43
16'b0000010000001110,        // LineF00 17.432at index 53
16'b0000010001000011,        // LineF00 18.333at index 60
16'b0000010001001101,        // LineF00 18.500at index 61
16'b0000010001011001,        // LineF00 18.698at index 62
16'b0000010100101001,        // LineF00 22.198at index 87
16'b0000010101011111,        // LineF00 23.099at index 93
16'b0000010101110011,        // LineF00 23.432at index 95
16'b0000010110001001,        // LineF00 23.798at index 98
16'b0000010110011100,        // LineF00 24.132at index 100
16'b0000010110110010,        // LineF00 24.499at index 103
16'b0000011001110001,        // LineF00 27.699at index 115
16'b0000011010000101,        // LineF00 28.032at index 117
16'b0000011010011010,        // LineF00 28.399at index 119
16'b0000011011100100,        // LineF00 29.632at index 125
16'b0000011100100011,        // LineF00 30.699at index 131
16'b0100011100110111,        // LineF01 31.031at index 133
16'b1000011101001101,        // LineF10 31.399at index 135
16'b0000011101101011,        // LineF00 31.898at index 139
16'b0000011110000011,        // LineF00 32.299at index 141
16'b0000011110010100,        // LineF00 32.584at index 144
16'b0000011110101100,        // LineF00 32.999at index 146
16'b0100100000110101,        // LineF01 35.300at index 160
16'b1000100001000111,        // LineF10 35.599at index 161
16'b0000100010001000,        // LineF00 36.698at index 166
16'b0000100010011100,        // LineF00 37.033at index 168
16'b0000100011011100,        // LineF00 38.098at index 179
16'b0100100011101000,        // LineF01 38.299at index 180
16'b1000100011110000,        // LineF10 38.431at index 182
16'b0000100100011001,        // LineF00 39.133at index 187
16'b0100100101000011,        // LineF01 39.832at index 195
16'b1000100101001111,        // LineF10 40.032at index 196
16'b0000100101111001,        // LineF00 40.734at index 201
16'b0000100111001100,        // LineF00 42.133at index 215
16'b0000100111110110,        // LineF00 42.833at index 221
16'b0100101000001011,        // LineF01 43.200at index 223
16'b1000101001111110,        // LineF10 45.133at index 233
16'b0000101010100000,        // LineF00 45.699at index 238
16'b0100101011101000,        // LineF01 46.898at index 245
16'b1000101011111111,        // LineF10 47.299at index 246
16'b0000101100011101,        // LineF00 47.798at index 250
16'b0000101100111101,        // LineF00 48.332at index 254
16'b0000101110010000,        // LineF00 49.731at index 261
16'b0000110000100011,        // LineF00 52.200at index 274
16'b0100110001001101,        // LineF01 52.899at index 279
16'b1000110001100101,        // LineF10 53.299at index 280
16'b0000110010010100,        // LineF00 54.099at index 285
16'b0100110011010110,        // LineF01 55.198at index 294
16'b1000110011101101,        // LineF10 55.599at index 295
16'b0000110100010001,        // LineF00 56.200at index 299
16'b0000110101101010,        // LineF00 57.699at index 308
16'b0000110110110010,        // LineF00 58.899at index 316
16'b0000111000010111,        // LineF00 60.598at index 322
16'b0000111010000100,        // LineF00 62.432at index 330
16'b0000111010011010,        // LineF00 62.798at index 334
16'b0000111010110100,        // LineF00 63.233at index 337
16'b0100111011011101,        // LineF01 63.932at index 340
16'b1000111100000111,        // LineF10 64.632at index 342
16'b0000111100011101,        // LineF00 65.000at index 344
16'b0000111100110101,        // LineF00 65.399at index 346
16'b0000111101011110,        // LineF00 66.098at index 350
16'b0000111110010000,        // LineF00 66.933at index 354
16'b0001000000011001,        // LineF00 69.233at index 368
16'b0001000001101100,        // LineF00 70.632at index 373
16'b0001000010111000,        // LineF00 71.899at index 382
16'b0001000011000100,        // LineF00 72.098at index 384
16'b0001000011010101,        // LineF00 72.398at index 388
16'b0001000100010111,        // LineF00 73.499at index 393
16'b0001000100110101,        // LineF00 73.998at index 395
16'b0101000101000001,        // LineF01 74.198at index 398
16'b1001000101010100,        // LineF10 74.532at index 399
16'b0001000101101010,        // LineF00 74.898at index 403
16'b0001000101111110,        // LineF00 75.233at index 407
16'b0001000110100100,        // LineF00 75.868at index 412
16'b0001000111001111,        // LineF00 76.599at index 415
16'b0001000111010111,        // LineF00 76.731at index 417
16'b0101000111100111,        // LineF01 76.999at index 420
16'b1001000111111111,        // LineF10 77.400at index 421
16'b0001001000011101,        // LineF00 77.899at index 424
16'b0001001001111100,        // LineF00 79.497at index 432
16'b0001001010001110,        // LineF00 79.798at index 434
16'b0001001010011010,        // LineF00 80.000at index 436
16'b0001001010100110,        // LineF00 80.199at index 438
16'b0001001100001101,        // LineF00 81.932at index 446
16'b0001001100011001,        // LineF00 82.133at index 448
16'b0001001101011100,        // LineF00 83.266at index 455
16'b0001001110011010,        // LineF00 84.300at index 463
16'b0001001111001101,        // LineF00 85.165at index 469
16'b0001001111100101,        // LineF00 85.566at index 471
16'b0001001111101101,        // LineF00 85.699at index 473
16'b0001001111110111,        // LineF00 85.865at index 474
16'b0001010001000001,        // LineF00 87.100at index 483
16'b0001010001101110,        // LineF00 87.867at index 488
16'b0001010011101011,        // LineF00 89.965at index 503
16'b0001010011110011,        // LineF00 90.098at index 505
16'b0001010011111101,        // LineF00 90.266at index 506
16'b0001010100001001,        // LineF00 90.466at index 507
16'b0001010101001010,        // LineF00 91.565at index 513
16'b0001010101110100,        // LineF00 92.265at index 518
16'b0001011001010011,
16'b0001011001010011,
16'b0001011001010011,
16'b0001011001010011
};

assign	key_1 = mem[addr];
assign	key_2 = mem[addr+1];
assign	key_3 = mem[addr+2];
assign	key_4 = mem[addr+3];

endmodule
