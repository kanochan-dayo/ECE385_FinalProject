module key_j(input [7:0] addr, 
output [15:0] key_1, 
output [15:0] key_2, 
output [15:0] key_3, 
output [15:0] key_4);
parameter [0:255][15:0] mem={
16'b0000000000110010,        // LineJ00 0.832at index 2
16'b0000000001010011,        // LineJ00 1.399at index 4
16'b0000000010110010,        // LineJ00 2.998at index 9
16'b0000000011011100,        // LineJ00 3.699at index 11
16'b0000000100000110,        // LineJ00 4.399at index 13
16'b0000000101000011,        // LineJ00 5.432at index 16
16'b0000000110100011,        // LineJ00 7.032at index 21
16'b0000000111001100,        // LineJ00 7.732at index 24
16'b0000001001010101,        // LineJ00 10.031at index 29
16'b0100001010101000,        // LineJ01 11.421at index 32
16'b1000001101010011,        // LineJ10 14.298at index 34
16'b0000001110111010,        // LineJ00 16.033at index 44
16'b0000001111000100,        // LineJ00 16.199at index 45
16'b0000001111010000,        // LineJ00 16.399at index 46
16'b0000001111011000,        // LineJ00 16.532at index 48
16'b0000010000000110,        // LineJ00 17.299at index 52
16'b0000010001100001,        // LineJ00 18.833at index 64
16'b0000010001101101,        // LineJ00 19.033at index 65
16'b0000010001110111,        // LineJ00 19.198at index 66
16'b0000010010000011,        // LineJ00 19.399at index 67
16'b0000010011000000,        // LineJ00 20.432at index 74
16'b0000010011101110,        // LineJ00 21.198at index 80
16'b0000010011110100,        // LineJ00 21.299at index 81
16'b0000010100000000,        // LineJ00 21.499at index 82
16'b0000010100001100,        // LineJ00 21.699at index 83
16'b0000010101101011,        // LineJ00 23.299at index 94
16'b0000010101111101,        // LineJ00 23.600at index 97
16'b0000010110010100,        // LineJ00 23.998at index 99
16'b0000010110101000,        // LineJ00 24.333at index 102
16'b0100010110111110,        // LineJ01 24.700at index 105
16'b1000011000011101,        // LineJ10 26.299at index 107
16'b0000011000100101,        // LineJ00 26.432at index 108
16'b0000011000111011,        // LineJ00 26.800at index 110
16'b0000011001001110,        // LineJ00 27.113at index 112
16'b0000011010111000,        // LineJ00 28.899at index 122
16'b0000011011100100,        // LineJ00 29.632at index 126
16'b0000011011111010,        // LineJ00 29.999at index 128
16'b0100011100001110,        // LineJ01 30.333at index 130
16'b1000011100100011,        // LineJ10 30.699at index 132
16'b0000011101001101,        // LineJ00 31.399at index 136
16'b0000011110000011,        // LineJ00 32.299at index 142
16'b0000011110101100,        // LineJ00 32.999at index 147
16'b0000011111001010,        // LineJ00 33.498at index 150
16'b0000011111110100,        // LineJ00 34.198at index 154
16'b0100100000001011,        // LineJ01 34.598at index 156
16'b1000100000011101,        // LineJ10 34.899at index 157
16'b0000100001110011,        // LineJ00 36.332at index 165
16'b0000100010001000,        // LineJ00 36.698at index 167
16'b0000100010110010,        // LineJ00 37.399at index 172
16'b0000100011000110,        // LineJ00 37.732at index 175
16'b0100100011110000,        // LineJ01 38.431at index 183
16'b1000100011111100,        // LineJ10 38.633at index 184
16'b0000100100101111,        // LineJ00 39.499at index 191
16'b0000100101011001,        // LineJ00 40.199at index 197
16'b0100100110011010,        // LineJ01 41.300at index 208
16'b1000100110100010,        // LineJ10 41.432at index 209
16'b0000100110111000,        // LineJ00 41.798at index 212
16'b0000101000000001,        // LineJ00 43.031at index 222
16'b0100101000110101,        // LineJ01 43.898at index 227
16'b1000101001000001,        // LineJ10 44.099at index 228
16'b0000101001110111,        // LineJ00 45.000at index 232
16'b0100101010101000,        // LineJ01 45.833at index 239
16'b1000101010111110,        // LineJ10 46.198at index 240
16'b0000101011011110,        // LineJ00 46.733at index 244
16'b0000101100010001,        // LineJ00 47.599at index 249
16'b0000101100110001,        // LineJ00 48.132at index 253
16'b0000101111101110,        // LineJ00 51.300at index 269
16'b0000110010010110,        // LineJ00 54.132at index 286
16'b0100110010101100,        // LineJ01 54.499at index 290
16'b1000110011000000,        // LineJ10 54.833at index 291
16'b0000110011111111,        // LineJ00 55.895at index 298
16'b0000110100010111,        // LineJ00 56.299at index 300
16'b0000110101011110,        // LineJ00 57.498at index 307
16'b0000110110001000,        // LineJ00 58.199at index 313
16'b0000110110110010,        // LineJ00 58.899at index 317
16'b0000110111111001,        // LineJ00 60.099at index 321
16'b0000111001000001,        // LineJ00 61.299at index 327
16'b0100111001110110,        // LineJ01 62.199at index 328
16'b1000111010000010,        // LineJ10 62.400at index 329
16'b0000111010010100,        // LineJ00 62.698at index 333
16'b0000111011001010,        // LineJ00 63.598at index 339
16'b0100111101000111,        // LineJ01 65.698at index 348
16'b1000111101011110,        // LineJ10 66.098at index 349
16'b0000111101111100,        // LineJ00 66.598at index 353
16'b0000111110100110,        // LineJ00 67.298at index 356
16'b0000111111000100,        // LineJ00 67.799at index 358
16'b0100111111101111,        // LineJ01 68.531at index 364
16'b1001000000000101,        // LineJ10 68.898at index 365
16'b0101000000101111,        // LineJ01 69.598at index 370
16'b1001000001011000,        // LineJ10 70.299at index 371
16'b0001000010001110,        // LineJ00 71.198at index 377
16'b0001000010101100,        // LineJ00 71.699at index 381
16'b0001000011000100,        // LineJ00 72.098at index 385
16'b0001000011001100,        // LineJ00 72.233at index 387
16'b0101000011100001,        // LineJ01 72.598at index 390
16'b1001000011111111,        // LineJ10 73.099at index 391
16'b0001000100110101,        // LineJ00 73.998at index 396
16'b0001000101011110,        // LineJ00 74.699at index 402
16'b0001000101101010,        // LineJ00 74.898at index 404
16'b0001000101111110,        // LineJ00 75.233at index 408
16'b0101000110001000,        // LineJ01 75.399at index 410
16'b1001000110100100,        // LineJ10 75.868at index 411
16'b0001000111001010,        // LineJ00 76.500at index 414
16'b0001000111111111,        // LineJ00 77.400at index 422
16'b0001001000110001,        // LineJ00 78.232at index 427
16'b0001001001010010,        // LineJ00 78.798at index 429
16'b0001001011000011,        // LineJ00 80.698at index 441
16'b0101001011011011,        // LineJ01 81.099at index 443
16'b1001001100000101,        // LineJ10 81.798at index 445
16'b0001001100010011,        // LineJ00 82.033at index 447
16'b0001001100011101,        // LineJ00 82.199at index 449
16'b0001001101111010,        // LineJ00 83.766at index 460
16'b0001001110011010,        // LineJ00 84.300at index 464
16'b0001001110100100,        // LineJ00 84.466at index 465
16'b0001001110110000,        // LineJ00 84.667at index 466
16'b0001010000000011,        // LineJ00 86.065at index 476
16'b0001010000001111,        // LineJ00 86.265at index 477
16'b0001010000010111,        // LineJ00 86.398at index 478
16'b0001010010001100,        // LineJ00 88.366at index 492
16'b0001010010011000,        // LineJ00 88.566at index 493
16'b0001010010100000,        // LineJ00 88.698at index 494
16'b0001010011001001,        // LineJ00 89.398at index 500
16'b0001010011010101,        // LineJ00 89.601at index 501
16'b0001010011011111,        // LineJ00 89.767at index 502
16'b0001010101010010,        // LineJ00 91.700at index 514
16'b0001010101101000,        // LineJ00 92.065at index 517
16'b0001011001010011,
16'b0001011001010011,
16'b0001011001010011,
16'b0001011001010011
};

assign	key_1 = mem[addr];
assign	key_2 = mem[addr+1];
assign	key_3 = mem[addr+2];
assign	key_4 = mem[addr+3];

endmodule
