module audio_clk_gen ();

endmodule