module arbiter ();

endmodule