module background_mapper (
);





endmodule