module frame_buffer(
input clk,
input [9:0] DrawX,     
				DrawY,
				ModX,     
				ModY,
				
input [3:0] MRed, MGreen, MBlue,
output logic [3:0]  Red, Green, Blue
);


endmodule