/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  background_palette_rom
(
		input [7:0] address,
		output logic [23:0] data_Out
);

// mem has width of 3 bits and a total of 400 addresses
parameter [0:255][23:0] mem ={

24'h000000,
24'h800000,
24'h008000,
24'h808000,
24'h000080,
24'h800080,
24'h008080,
24'hC0C0C0,
24'h808080,
24'hFF0000,
24'h00FF00,
24'hFFFF00,
24'h0000FF,
24'hFF00FF,
24'h00FFFF,
24'hFFFFFF,
24'h000000,
24'h00005F,
24'h000087,
24'h0000AF,
24'h0000D7,
24'h0000FF,
24'h005F00,
24'h005F5F,
24'h005F87,
24'h005FAF,
24'h005FD7,
24'h005FFF,
24'h008700,
24'h00875F,
24'h008787,
24'h0087AF,
24'h0087D7,
24'h0087FF,
24'h00AF00,
24'h00AF5F,
24'h00AF87,
24'h00AFAF,
24'h00AFD7,
24'h00AFFF,
24'h00D700,
24'h00D75F,
24'h00D787,
24'h00D7AF,
24'h00D7D7,
24'h00D7FF,
24'h00FF00,
24'h00FF5F,
24'h00FF87,
24'h00FFAF,
24'h00FFD7,
24'h00FFFF,
24'h5F0000,
24'h5F005F,
24'h5F0087,
24'h5F00AF,
24'h5F00D7,
24'h5F00FF,
24'h5F5F00,
24'h5F5F5F,
24'h5F5F87,
24'h5F5FAF,
24'h5F5FD7,
24'h5F5FFF,
24'h5F8700,
24'h5F875F,
24'h5F8787,
24'h5F87AF,
24'h5F87D7,
24'h5F87FF,
24'h5FAF00,
24'h5FAF5F,
24'h5FAF87,
24'h5FAFAF,
24'h5FAFD7,
24'h5FAFFF,
24'h5FD700,
24'h5FD75F,
24'h5FD787,
24'h5FD7AF,
24'h5FD7D7,
24'h5FD7FF,
24'h5FFF00,
24'h5FFF5F,
24'h5FFF87,
24'h5FFFAF,
24'h5FFFD7,
24'h5FFFFF,
24'h870000,
24'h87005F,
24'h870087,
24'h8700AF,
24'h8700D7,
24'h8700FF,
24'h875F00,
24'h875F5F,
24'h875F87,
24'h875FAF,
24'h875FD7,
24'h875FFF,
24'h878700,
24'h87875F,
24'h878787,
24'h8787AF,
24'h8787D7,
24'h8787FF,
24'h87AF00,
24'h87AF5F,
24'h87AF87,
24'h87AFAF,
24'h87AFD7,
24'h87AFFF,
24'h87D700,
24'h87D75F,
24'h87D787,
24'h87D7AF,
24'h87D7D7,
24'h87D7FF,
24'h87FF00,
24'h87FF5F,
24'h87FF87,
24'h87FFAF,
24'h87FFD7,
24'h87FFFF,
24'hAF0000,
24'hAF005F,
24'hAF0087,
24'hAF00AF,
24'hAF00D7,
24'hAF00FF,
24'hAF5F00,
24'hAF5F5F,
24'hAF5F87,
24'hAF5FAF,
24'hAF5FD7,
24'hAF5FFF,
24'hAF8700,
24'hAF875F,
24'hAF8787,
24'hAF87AF,
24'hAF87D7,
24'hAF87FF,
24'hAFAF00,
24'hAFAF5F,
24'hAFAF87,
24'hAFAFAF,
24'hAFAFD7,
24'hAFAFFF,
24'hAFD700,
24'hAFD75F,
24'hAFD787,
24'hAFD7AF,
24'hAFD7D7,
24'hAFD7FF,
24'hAFFF00,
24'hAFFF5F,
24'hAFFF87,
24'hAFFFAF,
24'hAFFFD7,
24'hAFFFFF,
24'hD70000,
24'hD7005F,
24'hD70087,
24'hD700AF,
24'hD700D7,
24'hD700FF,
24'hD75F00,
24'hD75F5F,
24'hD75F87,
24'hD75FAF,
24'hD75FD7,
24'hD75FFF,
24'hD78700,
24'hD7875F,
24'hD78787,
24'hD787AF,
24'hD787D7,
24'hD787FF,
24'hD7AF00,
24'hD7AF5F,
24'hD7AF87,
24'hD7AFAF,
24'hD7AFD7,
24'hD7AFFF,
24'hD7D700,
24'hD7D75F,
24'hD7D787,
24'hD7D7AF,
24'hD7D7D7,
24'hD7D7FF,
24'hD7FF00,
24'hD7FF5F,
24'hD7FF87,
24'hD7FFAF,
24'hD7FFD7,
24'hD7FFFF,
24'hFF0000,
24'hFF005F,
24'hFF0087,
24'hFF00AF,
24'hFF00D7,
24'hFF00FF,
24'hFF5F00,
24'hFF5F5F,
24'hFF5F87,
24'hFF5FAF,
24'hFF5FD7,
24'hFF5FFF,
24'hFF8700,
24'hFF875F,
24'hFF8787,
24'hFF87AF,
24'hFF87D7,
24'hFF87FF,
24'hFFAF00,
24'hFFAF5F,
24'hFFAF87,
24'hFFAFAF,
24'hFFAFD7,
24'hFFAFFF,
24'hFFD700,
24'hFFD75F,
24'hFFD787,
24'hFFD7AF,
24'hFFD7D7,
24'hFFD7FF,
24'hFFFF00,
24'hFFFF5F,
24'hFFFF87,
24'hFFFFAF,
24'hFFFFD7,
24'hFFFFFF,
24'h080808,
24'h121212,
24'h1C1C1C,
24'h262626,
24'h303030,
24'h3A3A3A,
24'h444444,
24'h4E4E4E,
24'h585858,
24'h626262,
24'h6C6C6C,
24'h767676,
24'h808080,
24'h8A8A8A,
24'h949494,
24'h9E9E9E,
24'hA8A8A8,
24'hB2B2B2,
24'hBCBCBC,
24'hC6C6C6,
24'hD0D0D0,
24'hDADADA,
24'hE4E4E4,
24'hEEEEEE
};


assign	data_Out = mem[address];


endmodule
