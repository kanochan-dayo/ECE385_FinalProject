//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//                                                                       --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 7                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------


module  color_mapper ( input        [9:0] DrawX, DrawY,
								input [31:0] data_in,
								input [11:0] fcolor_in,
								input [11:0] bcolor_in,
								input blank,
								input pixel_clk,
                       output logic [3:0]  Red, Green, Blue,
							 output logic[10:0] data_addr,
							 output logic[3:0] fcolor_addr,
							output logic[3:0] bcolor_addr	 );
    
	logic [10:0]	font_addr;
	logic [7:0]	font_data;
	logic num_of_char;
	logic [3:0] pix_row_of_char;
		
   font_rom ft_rom0(.addr(font_addr),.data(font_data));
	
	always_comb
	begin
	data_addr=DrawX[9:4]+DrawY[9:4]*40;
	pix_row_of_char=DrawY[3:0];
	num_of_char=DrawX[3];
	unique case(num_of_char)
	1'b0:
	begin
	font_addr={data_in[14:8],pix_row_of_char};
	fcolor_addr=data_in[7:4];
	bcolor_addr=data_in[3:0];
	end
	1'b1:
	begin
	font_addr={data_in[30:24],pix_row_of_char};
	fcolor_addr=data_in[23:20];
	bcolor_addr=data_in[19:16];
	end
	endcase
	end
	
	
	
	always_ff @(posedge pixel_clk)
	begin
	if(blank)
	case(font_data[7-DrawX[2:0]]^data_in[num_of_char*16+15])
	1'b1:
	begin
	Red<=fcolor_in[11:8];
	Green<=fcolor_in[7:4];
	Blue<=fcolor_in[3:0];
	end
	1'b0:
	begin
	Red<=bcolor_in[11:8];
	Green<=bcolor_in[7:4];
	Blue<=bcolor_in[3:0];
	end
	endcase
	else 
	begin
	Red<=0;
	Green<=0;
	Blue<=0;
	end
	end
	 
 /* Old Ball: Generated square box by checking if the current pixel is within a square of length
    2*Ball_Size, centered at (BallX, BallY).  Note that this requires unsigned comparisons.
	 
    if ((DrawX >= BallX - Ball_size) &&
       (DrawX <= BallX + Ball_size) &&
       (DrawY >= BallY - Ball_size) &&
       (DrawY <= BallY + Ball_size))

     New Ball: Generates (pixelated) circle by using the standard circle formula.  Note that while 
     this single line is quite powerful descriptively, it causes the synthesis tool to use up three
     of the 12 available multipliers on the chip!  Since the multiplicants are required to be signed,
	  we have to first cast them from logic to int (signed by default) before they are multiplied). */
	  
//    int DistX, DistY, Size;
//	 assign DistX = DrawX - BallX;
//    assign DistY = DrawY - BallY;
//    assign Size = Ball_size;
//	  
//    always_comb
//    begin:Ball_on_proc
//        if ( ( DistX*DistX + DistY*DistY) <= (Size * Size) ) 
//            ball_on = 1'b1;
//        else 
//            ball_on = 1'b0;
//     end 
//       
//    always_comb
//    begin:RGB_Display
//        if ((ball_on == 1'b1)) 
//        begin 
//            Red = 8'hff;
//            Green = 8'h55;
//            Blue = 8'h00;
//        end       
//        else 
//        begin 
//            Red = 8'h00; 
//            Green = 8'h00;
//            Blue = 8'h7f - DrawX[9:3];
//        end      
//    end 
    
endmodule
