module key_d(input [7:0] addr, 
output [15:0] key_1, 
output [15:0] key_2, 
output [15:0] key_3, 
output [15:0] key_4);
parameter [0:255][15:0] mem={
16'b0000000000110010,        \\ LineD00 0.832at index 1
16'b0000000011110000,        \\ LineD00 4.032at index 12
16'b0100000100011010,        \\ LineD01 4.731at index 14
16'b1000000101000011,        \\ LineD10 5.432at index 15
16'b0000000111001100,        \\ LineD00 7.732at index 23
16'b0000001000101010,        \\ LineD00 9.300at index 27
16'b0000001101111101,        \\ LineD00 14.999at index 35
16'b0000001110011011,        \\ LineD00 15.499at index 39
16'b0000001110100110,        \\ LineD00 15.698at index 41
16'b0000001110101110,        \\ LineD00 15.832at index 42
16'b0000001111011000,        \\ LineD00 16.532at index 47
16'b0000001111100100,        \\ LineD00 16.732at index 49
16'b0000001111101110,        \\ LineD00 16.898at index 50
16'b0000001111111010,        \\ LineD00 17.098at index 51
16'b0000010000100011,        \\ LineD00 17.799at index 55
16'b0000010001100001,        \\ LineD00 18.833at index 63
16'b0000010010000011,        \\ LineD00 19.399at index 68
16'b0000010010001111,        \\ LineD00 19.599at index 69
16'b0000010010010111,        \\ LineD00 19.732at index 70
16'b0000010010100000,        \\ LineD00 19.899at index 71
16'b0000010010111000,        \\ LineD00 20.298at index 73
16'b0000010011001010,        \\ LineD00 20.599at index 75
16'b0000010011010101,        \\ LineD00 20.783at index 77
16'b0000010011100010,        \\ LineD00 20.999at index 78
16'b0000010011101110,        \\ LineD00 21.198at index 79
16'b0000010100001100,        \\ LineD00 21.699at index 84
16'b0000010100010100,        \\ LineD00 21.833at index 85
16'b0000010100011111,        \\ LineD00 22.032at index 86
16'b0000010101111101,        \\ LineD00 23.600at index 96
16'b0000010110111110,        \\ LineD00 24.700at index 104
16'b0000011000011101,        \\ LineD00 26.299at index 106
16'b0000011000101111,        \\ LineD00 26.598at index 109
16'b0000011001000111,        \\ LineD00 26.999at index 111
16'b0000011001011001,        \\ LineD00 27.298at index 113
16'b0000011010101110,        \\ LineD00 28.733at index 121
16'b0000011011010000,        \\ LineD00 29.298at index 123
16'b0000011011111010,        \\ LineD00 29.999at index 127
16'b0000011100001110,        \\ LineD00 30.333at index 129
16'b0000011101011001,        \\ LineD00 31.599at index 137
16'b0000011111000000,        \\ LineD00 33.332at index 149
16'b0000011111010110,        \\ LineD00 33.701at index 151
16'b0000011111101010,        \\ LineD00 34.032at index 153
16'b0000100000000000,        \\ LineD00 34.400at index 155
16'b0000100000011101,        \\ LineD00 34.899at index 158
16'b0000100001011111,        \\ LineD00 35.998at index 163
16'b0000100010101100,        \\ LineD00 37.298at index 171
16'b0100100010111110,        \\ LineD01 37.600at index 173
16'b1000100011000110,        \\ LineD10 37.732at index 174
16'b0000100011010000,        \\ LineD00 37.898at index 176
16'b0100100100100011,        \\ LineD01 39.299at index 188
16'b1000100100101111,        \\ LineD10 39.499at index 190
16'b0000100100111011,        \\ LineD00 39.698at index 192
16'b0100100101011001,        \\ LineD01 40.199at index 198
16'b1000100101110001,        \\ LineD10 40.599at index 199
16'b0000100110000010,        \\ LineD00 40.899at index 204
16'b0100100110001110,        \\ LineD01 41.099at index 205
16'b1000100110011010,        \\ LineD10 41.300at index 207
16'b0100100110101100,        \\ LineD01 41.599at index 211
16'b1000100111000100,        \\ LineD10 41.998at index 213
16'b0100100111010110,        \\ LineD01 42.298at index 217
16'b1000100111101110,        \\ LineD10 42.699at index 219
16'b0000101010000100,        \\ LineD00 45.231at index 235
16'b0000101010010100,        \\ LineD00 45.499at index 237
16'b0000101010111110,        \\ LineD00 46.198at index 241
16'b0000101011010110,        \\ LineD00 46.598at index 243
16'b0000101100010001,        \\ LineD00 47.599at index 248
16'b0000101101000111,        \\ LineD00 48.499at index 255
16'b0000101101011011,        \\ LineD00 48.832at index 256
16'b0000101101110001,        \\ LineD00 49.199at index 259
16'b0100101110100110,        \\ LineD01 50.098at index 263
16'b1000101110111010,        \\ LineD10 50.431at index 265
16'b0000101111000100,        \\ LineD00 50.601at index 267
16'b0100101111111001,        \\ LineD01 51.499at index 270
16'b1000110000001101,        \\ LineD10 51.834at index 272
16'b0000110000111011,        \\ LineD00 52.599at index 277
16'b0000110001101101,        \\ LineD00 53.433at index 282
16'b0000110010000010,        \\ LineD00 53.799at index 283
16'b0000110010011100,        \\ LineD00 54.232at index 287
16'b0000110010101100,        \\ LineD00 54.499at index 289
16'b0000110011000000,        \\ LineD00 54.833at index 292
16'b0000110011111111,        \\ LineD00 55.895at index 297
16'b0100110100101001,        \\ LineD01 56.600at index 302
16'b1000110101000001,        \\ LineD10 56.998at index 303
16'b0000110101010101,        \\ LineD00 57.332at index 306
16'b0000110101110010,        \\ LineD00 57.833at index 310
16'b0000110110001000,        \\ LineD00 58.199at index 312
16'b0000110110100000,        \\ LineD00 58.599at index 314
16'b0000110110111110,        \\ LineD00 59.098at index 318
16'b0000110111111001,        \\ LineD00 60.099at index 320
16'b0000111000101011,        \\ LineD00 60.932at index 324
16'b0000111001000001,        \\ LineD00 61.299at index 326
16'b0000111010001110,        \\ LineD00 62.598at index 332
16'b0000111011001010,        \\ LineD00 63.598at index 338
16'b0000111101000111,        \\ LineD00 65.698at index 347
16'b0000111101111100,        \\ LineD00 66.598at index 352
16'b0000111110110010,        \\ LineD00 67.499at index 357
16'b0100111111000100,        \\ LineD01 67.799at index 359
16'b1000111111011011,        \\ LineD10 68.199at index 360
16'b0000111111100011,        \\ LineD00 68.333at index 362
16'b0000111111101111,        \\ LineD00 68.531at index 363
16'b0001000000000101,        \\ LineD00 68.898at index 366
16'b0001000000101111,        \\ LineD00 69.598at index 369
16'b0001000001011000,        \\ LineD00 70.299at index 372
16'b0001000010000010,        \\ LineD00 70.999at index 376
16'b0101000010010110,        \\ LineD01 71.332at index 379
16'b1001000010101100,        \\ LineD10 71.699at index 380
16'b0001000011001100,        \\ LineD00 72.233at index 386
16'b0001000011100001,        \\ LineD00 72.598at index 389
16'b0001000011111111,        \\ LineD00 73.099at index 392
16'b0001000101011110,        \\ LineD00 74.699at index 401
16'b0001000101110110,        \\ LineD00 75.098at index 405
16'b0001000110001000,        \\ LineD00 75.399at index 409
16'b0001000110111110,        \\ LineD00 76.299at index 413
16'b0001001000000111,        \\ LineD00 77.533at index 423
16'b0001001000110001,        \\ LineD00 78.232at index 426
16'b0001001001000110,        \\ LineD00 78.598at index 428
16'b0001001001100100,        \\ LineD00 79.098at index 430
16'b0001001010110010,        \\ LineD00 80.398at index 440
16'b0001001011011011,        \\ LineD00 81.099at index 442
16'b0001001011111001,        \\ LineD00 81.598at index 444
16'b0001001100100011,        \\ LineD00 82.298at index 450
16'b0001001100111011,        \\ LineD00 82.700at index 451
16'b0001001101000110,        \\ LineD00 82.899at index 453
16'b0001001101010000,        \\ LineD00 83.066at index 454
16'b0001001101111010,        \\ LineD00 83.766at index 459
16'b0001001110000110,        \\ LineD00 83.965at index 461
16'b0001001110001110,        \\ LineD00 84.107at index 462
16'b0001001110111000,        \\ LineD00 84.799at index 467
16'b0001010000000011,        \\ LineD00 86.065at index 475
16'b0001010000100001,        \\ LineD00 86.566at index 479
16'b0001010000101101,        \\ LineD00 86.765at index 481
16'b0001010000111001,        \\ LineD00 86.966at index 482
16'b0001010010000000,        \\ LineD00 88.165at index 490
16'b0001010010001100,        \\ LineD00 88.366at index 491
16'b0001010010101010,        \\ LineD00 88.866at index 495
16'b0001010010110110,        \\ LineD00 89.066at index 497
16'b0001010011000001,        \\ LineD00 89.265at index 498
16'b0001010011001001,        \\ LineD00 89.398at index 499
16'b0001010100011101,        \\ LineD00 90.799at index 509
16'b0001010100111110,        \\ LineD00 91.365at index 511
16'b0001010101011100,        \\ LineD00 91.865at index 515
16'b0101010101111100,        \\ LineD01 92.399at index 519
16'b1001010111100011,        \\ LineD10 94.133at index 521
};

assign	key_1 = mem[addr];
assign	key_2 = mem[addr+1];
assign	key_3 = mem[addr+2];
assign	key_4 = mem[addr+3];

endmodule
