module keycode_machine (
input [7:0] keycode,
input clk,reset,stop_sign,
output start_sign,
pause_sign,
result_ok
);

enum logic
endmodule
