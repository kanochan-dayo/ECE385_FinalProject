module arbiter_init(
input ram_init_done, 
);



endmodule