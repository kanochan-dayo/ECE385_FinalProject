/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  background_palette_rom
(
		input [7:0] address,
		output logic [23:0] data_Out
);

// mem has width of 3 bits and a total of 400 addresses
parameter [0:255][23:0] mem ={

24'h000000, 
24'h000050, 
24'h0000B0, 
24'h0000FF, 
24'h002000, 
24'h002050, 
24'h0020B0, 
24'h0020FF, 
24'h005000, 
24'h005050, 
24'h0050B0, 
24'h0050FF, 
24'h007000, 
24'h007050, 
24'h0070B0, 
24'h0070FF, 
24'h009000, 
24'h009050, 
24'h0090B0, 
24'h0090FF, 
24'h00B000, 
24'h00B050, 
24'h00B0B0, 
24'h00B0FF, 
24'h00E000, 
24'h00E050, 
24'h00E0B0, 
24'h00E0FF, 
24'h00FF00, 
24'h00FF50, 
24'h00FFB0, 
24'h00FFFF, 
24'h200000, 
24'h200050, 
24'h2000B0, 
24'h2000FF, 
24'h202000, 
24'h202050, 
24'h2020B0, 
24'h2020FF, 
24'h205000, 
24'h205050, 
24'h2050B0, 
24'h2050FF, 
24'h207000, 
24'h207050, 
24'h2070B0, 
24'h2070FF, 
24'h209000, 
24'h209050, 
24'h2090B0, 
24'h2090FF, 
24'h20B000, 
24'h20B050, 
24'h20B0B0, 
24'h20B0FF, 
24'h20E000, 
24'h20E050, 
24'h20E0B0, 
24'h20E0FF, 
24'h20FF00, 
24'h20FF50, 
24'h20FFB0, 
24'h20FFFF, 
24'h500000, 
24'h500050, 
24'h5000B0, 
24'h5000FF, 
24'h502000, 
24'h502050, 
24'h5020B0, 
24'h5020FF, 
24'h505000, 
24'h505050, 
24'h5050B0, 
24'h5050FF, 
24'h507000, 
24'h507050, 
24'h5070B0, 
24'h5070FF, 
24'h509000, 
24'h509050, 
24'h5090B0, 
24'h5090FF, 
24'h50B000, 
24'h50B050, 
24'h50B0B0, 
24'h50B0FF, 
24'h50E000, 
24'h50E050, 
24'h50E0B0, 
24'h50E0FF, 
24'h50FF00, 
24'h50FF50, 
24'h50FFB0, 
24'h50FFFF, 
24'h700000, 
24'h700050, 
24'h7000B0, 
24'h7000FF, 
24'h702000, 
24'h702050, 
24'h7020B0, 
24'h7020FF, 
24'h705000, 
24'h705050, 
24'h7050B0, 
24'h7050FF, 
24'h707000, 
24'h707050, 
24'h7070B0, 
24'h7070FF, 
24'h709000, 
24'h709050, 
24'h7090B0, 
24'h7090FF, 
24'h70B000, 
24'h70B050, 
24'h70B0B0, 
24'h70B0FF, 
24'h70E000, 
24'h70E050, 
24'h70E0B0, 
24'h70E0FF, 
24'h70FF00, 
24'h70FF50, 
24'h70FFB0, 
24'h70FFFF, 
24'h900000, 
24'h900050, 
24'h9000B0, 
24'h9000FF, 
24'h902000, 
24'h902050, 
24'h9020B0, 
24'h9020FF, 
24'h905000, 
24'h905050, 
24'h9050B0, 
24'h9050FF, 
24'h907000, 
24'h907050, 
24'h9070B0, 
24'h9070FF, 
24'h909000, 
24'h909050, 
24'h9090B0, 
24'h9090FF, 
24'h90B000, 
24'h90B050, 
24'h90B0B0, 
24'h90B0FF, 
24'h90E000, 
24'h90E050, 
24'h90E0B0, 
24'h90E0FF, 
24'h90FF00, 
24'h90FF50, 
24'h90FFB0, 
24'h90FFFF, 
24'hB00000, 
24'hB00050, 
24'hB000B0, 
24'hB000FF, 
24'hB02000, 
24'hB02050, 
24'hB020B0, 
24'hB020FF, 
24'hB05000, 
24'hB05050, 
24'hB050B0, 
24'hB050FF, 
24'hB07000, 
24'hB07050, 
24'hB070B0, 
24'hB070FF, 
24'hB09000, 
24'hB09050, 
24'hB090B0, 
24'hB090FF, 
24'hB0B000, 
24'hB0B050, 
24'hB0B0B0, 
24'hB0B0FF, 
24'hB0E000, 
24'hB0E050, 
24'hB0E0B0, 
24'hB0E0FF, 
24'hB0FF00, 
24'hB0FF50, 
24'hB0FFB0, 
24'hB0FFFF, 
24'hE00000, 
24'hE00050, 
24'hE000B0, 
24'hE000FF, 
24'hE02000, 
24'hE02050, 
24'hE020B0, 
24'hE020FF, 
24'hE05000, 
24'hE05050, 
24'hE050B0, 
24'hE050FF, 
24'hE07000, 
24'hE07050, 
24'hE070B0, 
24'hE070FF, 
24'hE09000, 
24'hE09050, 
24'hE090B0, 
24'hE090FF, 
24'hE0B000, 
24'hE0B050, 
24'hE0B0B0, 
24'hE0B0FF, 
24'hE0E000, 
24'hE0E050, 
24'hE0E0B0, 
24'hE0E0FF, 
24'hE0FF00, 
24'hE0FF50, 
24'hE0FFB0, 
24'hE0FFFF, 
24'hFF0000, 
24'hFF0050, 
24'hFF00B0, 
24'hFF00FF, 
24'hFF2000, 
24'hFF2050, 
24'hFF20B0, 
24'hFF20FF, 
24'hFF5000, 
24'hFF5050, 
24'hFF50B0, 
24'hFF50FF, 
24'hFF7000, 
24'hFF7050, 
24'hFF70B0, 
24'hFF70FF, 
24'hFF9000, 
24'hFF9050, 
24'hFF90B0, 
24'hFF90FF, 
24'hFFB000, 
24'hFFB050, 
24'hFFB0B0, 
24'hFFB0FF, 
24'hFFE000, 
24'hFFE050, 
24'hFFE0B0, 
24'hFFE0FF, 
24'hFFFF00, 
24'hFFFF50, 
24'hFFFFB0, 
24'hFFFFFF
};


assign	data_Out = mem[address];


endmodule
