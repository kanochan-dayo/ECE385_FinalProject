module key_k(input [7:0] addr, 
output [15:0] key_1, 
output [15:0] key_2, 
output [15:0] key_3, 
output [15:0] key_4
);
parameter [0:255][15:0] mem={
16'b0000000001100111,        // LineK00 1.732at index 5
16'b0000000001111101,        // LineK00 2.099at index 7
16'b0000000101011001,        // LineK00 5.799at index 17
16'b0000000110000011,        // LineK00 6.499at index 19
16'b0000001000011000,        // LineK00 8.998at index 26
16'b0000001001101011,        // LineK00 10.398at index 31
16'b0000001101111101,        // LineK00 14.999at index 36
16'b0000001110000101,        // LineK00 15.132at index 37
16'b0000001110001111,        // LineK00 15.299at index 38
16'b0000001110011011,        // LineK00 15.499at index 40
16'b0000010000011000,        // LineK00 17.599at index 54
16'b0000010000100011,        // LineK00 17.799at index 56
16'b0000010000101111,        // LineK00 18.000at index 57
16'b0000010000110111,        // LineK00 18.133at index 58
16'b0000010001000011,        // LineK00 18.333at index 59
16'b0000010010101100,        // LineK00 20.099at index 72
16'b0000010011001010,        // LineK00 20.599at index 76
16'b0000010100101001,        // LineK00 22.198at index 88
16'b0000010100110101,        // LineK00 22.398at index 89
16'b0000010100111101,        // LineK00 22.532at index 90
16'b0000010101001001,        // LineK00 22.733at index 91
16'b0000010101010011,        // LineK00 22.899at index 92
16'b0000010110011100,        // LineK00 24.132at index 101
16'b0000011001100101,        // LineK00 27.499at index 114
16'b0000011001111101,        // LineK00 27.898at index 116
16'b0000011010001111,        // LineK00 28.200at index 118
16'b0000011010100010,        // LineK00 28.532at index 120
16'b0000011011011000,        // LineK00 29.433at index 124
16'b0000011100110111,        // LineK00 31.031at index 134
16'b0000011101100001,        // LineK00 31.731at index 138
16'b0000011101110111,        // LineK00 32.101at index 140
16'b0000011110001011,        // LineK00 32.433at index 143
16'b0000011110100000,        // LineK00 32.800at index 145
16'b0000011110110100,        // LineK00 33.131at index 148
16'b0000011111011110,        // LineK00 33.833at index 152
16'b0000100000101001,        // LineK00 35.099at index 159
16'b0000100001000111,        // LineK00 35.599at index 162
16'b0000100001011111,        // LineK00 35.998at index 164
16'b0000100010011100,        // LineK00 37.033at index 169
16'b0000100010100110,        // LineK00 37.199at index 170
16'b0100100011010000,        // LineK01 37.898at index 177
16'b1000100011011100,        // LineK10 38.098at index 178
16'b0000100011101000,        // LineK00 38.299at index 181
16'b0100100100000101,        // LineK01 38.799at index 185
16'b1000100100011001,        // LineK10 39.133at index 186
16'b0000100100100011,        // LineK00 39.299at index 189
16'b0100100100111011,        // LineK01 39.698at index 193
16'b1000100101000011,        // LineK10 39.832at index 194
16'b0000100101110001,        // LineK00 40.599at index 200
16'b0100100101111001,        // LineK01 40.734at index 202
16'b1000100110000010,        // LineK10 40.899at index 203
16'b0000100110001110,        // LineK00 41.099at index 206
16'b0000100110101100,        // LineK00 41.599at index 210
16'b0100100111000100,        // LineK01 41.998at index 214
16'b1000100111010110,        // LineK10 42.298at index 216
16'b0000100111100010,        // LineK00 42.498at index 218
16'b0000100111101110,        // LineK00 42.699at index 220
16'b0100101000001011,        // LineK01 43.200at index 224
16'b1000101000010111,        // LineK10 43.398at index 225
16'b0000101000100011,        // LineK00 43.599at index 226
16'b0000101001001101,        // LineK00 44.300at index 229
16'b0100101001011111,        // LineK01 44.600at index 230
16'b1000101001101011,        // LineK10 44.798at index 231
16'b0000101001111110,        // LineK00 45.133at index 234
16'b0000101010001000,        // LineK00 45.299at index 236
16'b0000101011001010,        // LineK00 46.398at index 242
16'b0000101011111111,        // LineK00 47.299at index 247
16'b0000101100011101,        // LineK00 47.798at index 251
16'b0000101100101001,        // LineK00 48.000at index 252
16'b0100101101011011,        // LineK01 48.832at index 257
16'b1000101101110001,        // LineK10 49.199at index 258
16'b0000101101111100,        // LineK00 49.398at index 260
16'b0000101110010000,        // LineK00 49.731at index 262
16'b0000101110100110,        // LineK00 50.098at index 264
16'b0000101110111010,        // LineK00 50.431at index 266
16'b0000101111011100,        // LineK00 50.999at index 268
16'b0000101111111001,        // LineK00 51.499at index 271
16'b0000110000001101,        // LineK00 51.834at index 273
16'b0100110000100011,        // LineK01 52.200at index 275
16'b1000110000111011,        // LineK10 52.599at index 276
16'b0000110001001101,        // LineK00 52.899at index 278
16'b0000110001100101,        // LineK00 53.299at index 281
16'b0000110010001110,        // LineK00 53.999at index 284
16'b0000110010100000,        // LineK00 54.298at index 288
16'b0000110011010110,        // LineK00 55.198at index 293
16'b0000110011101101,        // LineK00 55.599at index 296
16'b0000110100101001,        // LineK00 56.600at index 301
16'b0100110101000001,        // LineK01 56.998at index 304
16'b1000110101010101,        // LineK10 57.332at index 305
16'b0000110101101010,        // LineK00 57.699at index 309
16'b0000110101110010,        // LineK00 57.833at index 311
16'b0000110110100000,        // LineK00 58.599at index 315
16'b0000110110111110,        // LineK00 59.098at index 319
16'b0000111000010111,        // LineK00 60.598at index 323
16'b0000111000101011,        // LineK00 60.932at index 325
16'b0000111010001010,        // LineK00 62.532at index 331
16'b0100111010100000,        // LineK01 62.898at index 335
16'b1000111010110100,        // LineK10 63.233at index 336
16'b0100111011011101,        // LineK01 63.932at index 341
16'b1000111100000111,        // LineK10 64.632at index 343
16'b0000111100011101,        // LineK00 65.000at index 345
16'b0000111101100110,        // LineK00 66.232at index 351
16'b0000111110010000,        // LineK00 66.933at index 355
16'b0000111111011011,        // LineK00 68.199at index 361
16'b0001000000011001,        // LineK00 69.233at index 367
16'b0001000001101100,        // LineK00 70.632at index 374
16'b0001000001111000,        // LineK00 70.833at index 375
16'b0001000010010110,        // LineK00 71.332at index 378
16'b0001000010111000,        // LineK00 71.899at index 383
16'b0001000100101000,        // LineK00 73.778at index 394
16'b0001000101000001,        // LineK00 74.198at index 397
16'b0001000101010100,        // LineK00 74.532at index 400
16'b0001000101110110,        // LineK00 75.098at index 406
16'b0001000111010001,        // LineK00 76.633at index 416
16'b0001000111011011,        // LineK00 76.797at index 418
16'b0001000111100111,        // LineK00 76.999at index 419
16'b0001001000011101,        // LineK00 77.899at index 425
16'b0001001001100100,        // LineK00 79.098at index 431
16'b0001001001111100,        // LineK00 79.497at index 433
16'b0001001010001110,        // LineK00 79.798at index 435
16'b0001001010011010,        // LineK00 80.000at index 437
16'b0001001010100110,        // LineK00 80.199at index 439
16'b0001001100111011,        // LineK00 82.700at index 452
16'b0001001101011100,        // LineK00 83.266at index 456
16'b0001001101100100,        // LineK00 83.398at index 457
16'b0001001101110000,        // LineK00 83.600at index 458
16'b0001001111000011,        // LineK00 84.999at index 468
16'b0001001111011001,        // LineK00 85.365at index 470
16'b0001001111100101,        // LineK00 85.566at index 472
16'b0001010000100001,        // LineK00 86.566at index 480
16'b0001010001000001,        // LineK00 87.100at index 484
16'b0001010001001100,        // LineK00 87.298at index 485
16'b0001010001010110,        // LineK00 87.465at index 486
16'b0001010001100010,        // LineK00 87.666at index 487
16'b0001010001110110,        // LineK00 87.998at index 489
16'b0001010010101010,        // LineK00 88.866at index 496
16'b0001010011101011,        // LineK00 89.965at index 504
16'b0001010100010101,        // LineK00 90.665at index 508
16'b0001010100101001,        // LineK00 90.999at index 510
16'b0001010100111110,        // LineK00 91.365at index 512
16'b0001010101011100,        // LineK00 91.865at index 516
16'b0101010101111100,        // LineK01 92.399at index 520
16'b1001010111100011,       // LineK10 94.133at index 522
16'b0001011001010011,
16'b0001011001010011,
16'b0001011001010011,
16'b0001011001010011,
};

assign	key_1 = mem[addr];
assign	key_2 = mem[addr+1];
assign	key_3 = mem[addr+2];
assign	key_4 = mem[addr+3];

endmodule
